module HALFSUB_BEHAV
(
input a,b,
output Borr,Diff
);

assign{Borr,Diff}=a-b;
endmodule
