module HA_BEHAV
(
input a,b,
output sum,Cout
);

assign{Cout,sum}=a+b;
endmodule
