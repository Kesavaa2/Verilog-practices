module pari_gen_odd
  (input a,b,c,
   output p);
  
  wire x;
      
  xor r1(x,b,c);
  xor r2(p,x,a);
endmodule
