module FA_BEHAV
(
input a,b,c,
output sum,Cout
);

assign{Cout,sum}=a+b+c;
endmodule
